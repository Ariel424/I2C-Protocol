//==============================================================================
// Testbench Top Module
//==============================================================================
module tb;
    
    //--------------------------------------------------------------------------
    // Testbench Components
    //--------------------------------------------------------------------------
    generator   gen;
    driver      drv;
    monitor     mon;
    scoreboard  sco;
    
    //--------------------------------------------------------------------------
    // Events
    //--------------------------------------------------------------------------
    event nextgd;
    event nextgs;
    
    //--------------------------------------------------------------------------
    // Mailboxes
    //--------------------------------------------------------------------------
    mailbox #(transaction) mbxgd, mbxms;
    
    //--------------------------------------------------------------------------
    // Interface and DUT Instantiation
    //--------------------------------------------------------------------------
    i2c_if vif();
    
    i2c_top dut (
        .clk     (vif.clk),
        .rst     (vif.rst),
        .newd    (vif.newd),
        .op      (vif.op),
        .addr    (vif.addr),
        .din     (vif.din),
        .dout    (vif.dout),
        .busy    (vif.busy),
        .ack_err (vif.ack_err),
        .done    (vif.done)
    );
    
    //--------------------------------------------------------------------------
    // Clock Generation
    //--------------------------------------------------------------------------
    initial begin
        vif.clk <= 0;
    end
    
    always #5 vif.clk <= ~vif.clk;
    
    //--------------------------------------------------------------------------
    // Testbench Initialization
    //--------------------------------------------------------------------------
    initial begin
        // Create mailboxes
        mbxgd = new();
        mbxms = new();
        
        // Create testbench components
        gen = new(mbxgd);
        drv = new(mbxgd);
        mon = new(mbxms);
        sco = new(mbxms);
        
        // Configure generator
        gen.count = 20;
        
        // Connect interfaces
        drv.vif = vif;
        mon.vif = vif;
        
        // Connect events
        gen.drvnext = nextgd;
        drv.drvnext = nextgd;
        gen.sconext = nextgs;
        sco.sconext = nextgs;
    end
    
    //--------------------------------------------------------------------------
    // Pre-Test Task
    //--------------------------------------------------------------------------
    task pre_test;
        drv.reset();
    endtask
    
    //--------------------------------------------------------------------------
    // Test Task
    //--------------------------------------------------------------------------
    task test;
        fork
            gen.run();
            drv.run();
            mon.run();
            sco.run();
        join_any
    endtask
    
    //--------------------------------------------------------------------------
    // Post-Test Task
    //--------------------------------------------------------------------------
    task post_test;
        wait(gen.done.triggered);
        $finish();
    endtask
    
    //--------------------------------------------------------------------------
    // Run Task
    //--------------------------------------------------------------------------
    task run();
        pre_test;
        test;
        post_test;
    endtask
    
    //--------------------------------------------------------------------------
    // Main Test Execution
    //--------------------------------------------------------------------------
    initial begin
        run();
    end
    
    //--------------------------------------------------------------------------
    // Waveform Dump
    //--------------------------------------------------------------------------
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars();
    end
    
endmodule
